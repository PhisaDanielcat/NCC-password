`timescale 1ns / 1ps

module S_box(
    input [7:0] inbox,
    output reg[7:0] outbox
    );
    
    always@(*)begin
        case(inbox)
            8'h00:outbox = 8'hd6;
            8'h01:outbox = 8'h90;
            8'h02:outbox = 8'he9;
            8'h03:outbox = 8'hfe;
            8'h04:outbox = 8'hcc;
            8'h05:outbox = 8'he1;
            8'h06:outbox = 8'h3d;
            8'h07:outbox = 8'hb7;
            8'h08:outbox = 8'h16;
            8'h09:outbox = 8'hb6;
            8'h0a:outbox = 8'h14;
            8'h0b:outbox = 8'hc2;
            8'h0c:outbox = 8'h28;
            8'h0d:outbox = 8'hfb;
            8'h0e:outbox = 8'h2c;
            8'h0f:outbox = 8'h05;
            8'h10:outbox = 8'h2b;
            8'h11:outbox = 8'h67;
            8'h12:outbox = 8'h9a;
            8'h13:outbox = 8'h76;
            8'h14:outbox = 8'h2a;
            8'h15:outbox = 8'hbe;
            8'h16:outbox = 8'h04;
            8'h17:outbox = 8'hc3;
            8'h18:outbox = 8'haa;
            8'h19:outbox = 8'h44;
            8'h1a:outbox = 8'h13;
            8'h1b:outbox = 8'h26;
            8'h1c:outbox = 8'h49;
            8'h1d:outbox = 8'h86;
            8'h1e:outbox = 8'h06;
            8'h1f:outbox = 8'h99;
            8'h20:outbox = 8'h9c;
            8'h21:outbox = 8'h42;
            8'h22:outbox = 8'h50;
            8'h23:outbox = 8'hf4;
            8'h24:outbox = 8'h91;
            8'h25:outbox = 8'hef;
            8'h26:outbox = 8'h98;
            8'h27:outbox = 8'h7a;
            8'h28:outbox = 8'h33;
            8'h29:outbox = 8'h54;
            8'h2a:outbox = 8'h0b;
            8'h2b:outbox = 8'h43;
            8'h2c:outbox = 8'hed;
            8'h2d:outbox = 8'hcf;
            8'h2e:outbox = 8'hac;
            8'h2f:outbox = 8'h62;
            8'h30:outbox = 8'he4;
            8'h31:outbox = 8'hb3;
            8'h32:outbox = 8'h1c;
            8'h33:outbox = 8'ha9;
            8'h34:outbox = 8'hc9;
            8'h35:outbox = 8'h08;
            8'h36:outbox = 8'he8;
            8'h37:outbox = 8'h95;
            8'h38:outbox = 8'h80;
            8'h39:outbox = 8'hdf;
            8'h3a:outbox = 8'h94;
            8'h3b:outbox = 8'hfa;
            8'h3c:outbox = 8'h75;
            8'h3d:outbox = 8'h8f;
            8'h3e:outbox = 8'h3f;
            8'h3f:outbox = 8'ha6;
            8'h40:outbox = 8'h47;
            8'h41:outbox = 8'h07;
            8'h42:outbox = 8'ha7;
            8'h43:outbox = 8'hfc;
            8'h44:outbox = 8'hf3;
            8'h45:outbox = 8'h73;
            8'h46:outbox = 8'h17;
            8'h47:outbox = 8'hba;
            8'h48:outbox = 8'h83;
            8'h49:outbox = 8'h59;
            8'h4a:outbox = 8'h3c;
            8'h4b:outbox = 8'h19;
            8'h4c:outbox = 8'he6;
            8'h4d:outbox = 8'h85;
            8'h4e:outbox = 8'h4f;
            8'h4f:outbox = 8'ha8;
            8'h50:outbox = 8'h68;
            8'h51:outbox = 8'h6b;
            8'h52:outbox = 8'h81;
            8'h53:outbox = 8'hb2;
            8'h54:outbox = 8'h71;
            8'h55:outbox = 8'h64;
            8'h56:outbox = 8'hda;
            8'h57:outbox = 8'h8b;
            8'h58:outbox = 8'hf8;
            8'h59:outbox = 8'heb;
            8'h5a:outbox = 8'h0f;
            8'h5b:outbox = 8'h4b;
            8'h5c:outbox = 8'h70;
            8'h5d:outbox = 8'h56;
            8'h5e:outbox = 8'h9d;
            8'h5f:outbox = 8'h35;
            8'h60:outbox = 8'h1e;
            8'h61:outbox = 8'h24;
            8'h62:outbox = 8'h0e;
            8'h63:outbox = 8'h5e;
            8'h64:outbox = 8'h63;
            8'h65:outbox = 8'h58;
            8'h66:outbox = 8'hd1;
            8'h67:outbox = 8'ha2;
            8'h68:outbox = 8'h25;
            8'h69:outbox = 8'h22;
            8'h6a:outbox = 8'h7c;
            8'h6b:outbox = 8'h3b;
            8'h6c:outbox = 8'h01;
            8'h6d:outbox = 8'h21;
            8'h6e:outbox = 8'h78;
            8'h6f:outbox = 8'h87;
            8'h70:outbox = 8'hd4;
            8'h71:outbox = 8'h00;
            8'h72:outbox = 8'h46;
            8'h73:outbox = 8'h57;
            8'h74:outbox = 8'h9f;
            8'h75:outbox = 8'hd3;
            8'h76:outbox = 8'h27;
            8'h77:outbox = 8'h52;
            8'h78:outbox = 8'h4c;
            8'h79:outbox = 8'h36;
            8'h7a:outbox = 8'h02;
            8'h7b:outbox = 8'he7;
            8'h7c:outbox = 8'ha0;
            8'h7d:outbox = 8'hc4;
            8'h7e:outbox = 8'hc8;
            8'h7f:outbox = 8'h9e;
            8'h80:outbox = 8'hea;
            8'h81:outbox = 8'hbf;
            8'h82:outbox = 8'h8a;
            8'h83:outbox = 8'hd2;
            8'h84:outbox = 8'h40;
            8'h85:outbox = 8'hc7;
            8'h86:outbox = 8'h38;
            8'h87:outbox = 8'hb5;
            8'h88:outbox = 8'ha3;
            8'h89:outbox = 8'hf7;
            8'h8a:outbox = 8'hf2;
            8'h8b:outbox = 8'hce;
            8'h8c:outbox = 8'hf9;
            8'h8d:outbox = 8'h61;
            8'h8e:outbox = 8'h15;
            8'h8f:outbox = 8'ha1;
            8'h90:outbox = 8'he0;
            8'h91:outbox = 8'hae;
            8'h92:outbox = 8'h5d;
            8'h93:outbox = 8'ha4;
            8'h94:outbox = 8'h9b;
            8'h95:outbox = 8'h34;
            8'h96:outbox = 8'h1a;
            8'h97:outbox = 8'h55;
            8'h98:outbox = 8'had;
            8'h99:outbox = 8'h93;
            8'h9a:outbox = 8'h32;
            8'h9b:outbox = 8'h30;
            8'h9c:outbox = 8'hf5;
            8'h9d:outbox = 8'h8c;
            8'h9e:outbox = 8'hb1;
            8'h9f:outbox = 8'he3;
            8'ha0:outbox = 8'h1d;
            8'ha1:outbox = 8'hf6;
            8'ha2:outbox = 8'he2;
            8'ha3:outbox = 8'h2e;
            8'ha4:outbox = 8'h82;
            8'ha5:outbox = 8'h66;
            8'ha6:outbox = 8'hca;
            8'ha7:outbox = 8'h60;
            8'ha8:outbox = 8'hc0;
            8'ha9:outbox = 8'h29;
            8'haa:outbox = 8'h23;
            8'hab:outbox = 8'hab;
            8'hac:outbox = 8'h0d;
            8'had:outbox = 8'h53;
            8'hae:outbox = 8'h4e;
            8'haf:outbox = 8'h6f;
            8'hb0:outbox = 8'hd5;
            8'hb1:outbox = 8'hdb;
            8'hb2:outbox = 8'h37;
            8'hb3:outbox = 8'h45;
            8'hb4:outbox = 8'hde;
            8'hb5:outbox = 8'hfd;
            8'hb6:outbox = 8'h8e;
            8'hb7:outbox = 8'h2f;
            8'hb8:outbox = 8'h03;
            8'hb9:outbox = 8'hff;
            8'hba:outbox = 8'h6a;
            8'hbb:outbox = 8'h72;
            8'hbc:outbox = 8'h6d;
            8'hbd:outbox = 8'h6c;
            8'hbe:outbox = 8'h5b;
            8'hbf:outbox = 8'h51;
            8'hc0:outbox = 8'h8d;
            8'hc1:outbox = 8'h1b;
            8'hc2:outbox = 8'haf;
            8'hc3:outbox = 8'h92;
            8'hc4:outbox = 8'hbb;
            8'hc5:outbox = 8'hdd;
            8'hc6:outbox = 8'hbc;
            8'hc7:outbox = 8'h7f;
            8'hc8:outbox = 8'h11;
            8'hc9:outbox = 8'hd9;
            8'hca:outbox = 8'h5c;
            8'hcb:outbox = 8'h41;
            8'hcc:outbox = 8'h1f;
            8'hcd:outbox = 8'h10;
            8'hce:outbox = 8'h5a;
            8'hcf:outbox = 8'hd8;
            8'hd0:outbox = 8'h0a;
            8'hd1:outbox = 8'hc1;
            8'hd2:outbox = 8'h31;
            8'hd3:outbox = 8'h88;
            8'hd4:outbox = 8'ha5;
            8'hd5:outbox = 8'hcd;
            8'hd6:outbox = 8'h7b;
            8'hd7:outbox = 8'hbd;
            8'hd8:outbox = 8'h2d;
            8'hd9:outbox = 8'h74;
            8'hda:outbox = 8'hd0;
            8'hdb:outbox = 8'h12;
            8'hdc:outbox = 8'hb8;
            8'hdd:outbox = 8'he5;
            8'hde:outbox = 8'hb4;
            8'hdf:outbox = 8'hb0;
            8'he0:outbox = 8'h89;
            8'he1:outbox = 8'h69;
            8'he2:outbox = 8'h97;
            8'he3:outbox = 8'h4a;
            8'he4:outbox = 8'h0c;
            8'he5:outbox = 8'h96;
            8'he6:outbox = 8'h77;
            8'he7:outbox = 8'h7e;
            8'he8:outbox = 8'h65;
            8'he9:outbox = 8'hb9;
            8'hea:outbox = 8'hf1;
            8'heb:outbox = 8'h09;
            8'hec:outbox = 8'hc5;
            8'hed:outbox = 8'h6e;
            8'hee:outbox = 8'hc6;
            8'hef:outbox = 8'h84;
            8'hf0:outbox = 8'h18;
            8'hf1:outbox = 8'hf0;
            8'hf2:outbox = 8'h7d;
            8'hf3:outbox = 8'hec;
            8'hf4:outbox = 8'h3a;
            8'hf5:outbox = 8'hdc;
            8'hf6:outbox = 8'h4d;
            8'hf7:outbox = 8'h20;
            8'hf8:outbox = 8'h79;
            8'hf9:outbox = 8'hee;
            8'hfa:outbox = 8'h5f;
            8'hfb:outbox = 8'h3e;
            8'hfc:outbox = 8'hd7;
            8'hfd:outbox = 8'hcb;
            8'hfe:outbox = 8'h39;
            8'hff:outbox = 8'h48;
        endcase
    end
endmodule
